package elevator_pkg;
   typedef enum reg {UP, DOWN} Direction;
   typedef enum reg {OPEN, CLOSE} DoorsOp;
   typedef enum reg {GO, STOP} EngineOp;
endpackage // elevator_pkg

